/*
 * Copyright (c) 2024 Fabio Ramirez Stern
 * SPDX-License-Identifier: Apache-2.0
 */

`define default_netname none

module tt_um_faramire_gate_guesser (
    input  wire [7:0] ui_in,    // Dedicated inputs:   switches 0 to 7
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path:    switches 8 to F
    output wire [7:0] uio_out,  // IOs: Output path:   gate outputs
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // will go high when the design is enabled
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // All output pins must be assigned. If not used, assign to 0.

    //TODO

  assign uo_out  = 0;
  assign uio_out = 0;
  assign uio_oe  = 0;

endmodule
